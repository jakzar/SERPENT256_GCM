library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.env.stop;

entity tb_serpent_dec is
end tb_serpent_dec;

architecture behavior of tb_serpent_dec is

    constant inClkp : time := 10ns;
    signal in_clk : std_logic := '0';

    signal in_reset : std_logic := '0';
    signal in_data      :  std_logic_vector (127 downto 0);
    signal in_key      :  std_logic_vector (255 downto 0);
    signal out_data      :  std_logic_vector (127 downto 0);

    signal in_key_wr  : std_logic;
    signal in_data_wr  : std_logic;

    signal out_busy  : std_logic;

begin
    in_clk <= not in_clk after inClkp/2;
    uut: entity work.serpent_dec port map(in_clk, in_reset, in_key_wr, in_data_wr, in_data, in_key, out_data, out_busy);
    process
        
    begin
        wait for 10 ns;
        wait for 10 ns;
        in_key_wr <= '1';
        in_data_wr <= '1';
        in_key<=x"3F9EE37D9EA55DAA6AB3911773F9C3E3EE74FED44397F0B6CF202CA0FE0903B7";
        in_data<=x"2868B7A2D28ECD5E4FDEFAC3C4330074";

        wait for 10 ns;
        in_key_wr <= '0';
        in_data_wr <= '0';
        in_key <= (others => '0');
        in_data <= (others => '0');
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        in_key_wr <= '1';
        in_data_wr <= '1';
        in_key<=x"8BF47F58C4A0518E2FE30405C4B637F9B465955B7D1F0BA7455BFD0739E3A810";
        in_data<=x"6AC7579D9377845A816CA6D758F3FEFF";
        wait for 10 ns;
        in_key_wr <= '0';
        in_data_wr <= '0';
        in_key <= (others => '0');
        in_data <= (others => '0');
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        in_key_wr <= '1';
        in_data_wr <= '1';
        in_key<=x"3F9EE37D9EA55DAA6AB3911773F9C3E3EE74FED44397F0B6CF202CA0FE0903B7";
        in_data<=x"2868B7A2D28ECD5E4FDEFAC3C4330074";

        wait for 10 ns;
        in_key_wr <= '0';
        in_data_wr <= '0';
        in_key <= (others => '0');
        in_data <= (others => '0');
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        in_reset<='1';
        wait for 10 ns;
        in_reset<='0';
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        in_key_wr <= '1';
        in_data_wr <= '1';
        in_key<=x"3F9EE37D9EA55DAA6AB3911773F9C3E3EE74FED44397F0B6CF202CA0FE0903B7";
        in_data<=x"2868B7A2D28ECD5E4FDEFAC3C4330074";

        wait for 10 ns;
        in_key_wr <= '0';
        in_data_wr <= '0';
        in_key <= (others => '0');
        in_data <= (others => '0');
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        wait for 10 ns;
        stop;
    end process;

end behavior;
